package Packet;

  class Packet;
    int field1; 

    function new(int i);
      field1 = i;
    endfunction   
  endclass : Packet

endpackage